//
//
//
//
//
//
//
//
`timescale 1ns / 1ps

//
module const0(out);
//
output [0:0] out;

//
//


//
//

	assign out[0] = 1'b0;
endmodule
//

//
module const1(const1);
//
output [0:0] const1;

//
//


//
//

	assign const1[0] = 1'b1;
endmodule
//

